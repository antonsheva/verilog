//====================================================================================================================================
module frFilter(
	CLK50, IN, OUT
);
	
	parameter MAX_CNT = 2'h1;
	parameter CNT_WIDTH = 2'h2;

	input CLK50, IN;
	output reg OUT;

//====================================================================================================================================

reg [(CNT_WIDTH-1):0] cnt;

always @(posedge CLK50) begin
	if(IN==OUT) cnt <= MAX_CNT;
	else begin
		if(cnt) cnt <= cnt - 1'b1;
		else begin
			OUT <= ~OUT;
			cnt <= MAX_CNT;
		end
	end
end

//====================================================================================================================================

endmodule
